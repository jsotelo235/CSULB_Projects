`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:17:11 04/23/2017 
// Design Name: 
// Module Name:    ram_1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ram_1(
    input clk,
    input we,
    input [15:0] addr,
    input [15:0] din,
    output [15:0] dout
    );


endmodule
